module invert(A, A_inv);
        
    input [31:0] A;
    output [31:0] A_inv;

    not not1(A_inv[0], A[0]);
    not not2(A_inv[1], A[1]);
    not not3(A_inv[2], A[2]);
    not not4(A_inv[3], A[3]);
    not not5(A_inv[4], A[4]);
    not not6(A_inv[5], A[5]);
    not not7(A_inv[6], A[6]);
    not not8(A_inv[7], A[7]);
    not not9(A_inv[8], A[8]);
    not not10(A_inv[9], A[9]);
    not not11(A_inv[10], A[10]);
    not not12(A_inv[11], A[11]);
    not not13(A_inv[12], A[12]);
    not not14(A_inv[13], A[13]);
    not not15(A_inv[14], A[14]);
    not not16(A_inv[15], A[15]);
    not not17(A_inv[16], A[16]);
    not not18(A_inv[17], A[17]);
    not not19(A_inv[18], A[18]);
    not not20(A_inv[19], A[19]);
    not not21(A_inv[20], A[20]);
    not not22(A_inv[21], A[21]);
    not not23(A_inv[22], A[22]);
    not not24(A_inv[23], A[23]);
    not not25(A_inv[24], A[24]);
    not not26(A_inv[25], A[25]);
    not not27(A_inv[26], A[26]);
    not not28(A_inv[27], A[27]);
    not not29(A_inv[28], A[28]);
    not not30(A_inv[29], A[29]);
    not not31(A_inv[30], A[30]);
    not not32(A_inv[31], A[31]);

endmodule